CircuitMaker Text
5.6
Probes: 1
Is2_1
Transient Analysis
0 415 44 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
347 79 1918 443
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.603191 0.500000
515 175 2086 742
9961490 0
0
6 Title:
5 Name:
0
0
0
27
7 Ground~
168 714 100 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3623 0 0
2
5.8993e-315 0
0
7 Ground~
168 755 102 0 1 3
0 2
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3722 0 0
2
5.8993e-315 5.38788e-315
0
7 Ground~
168 651 102 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8993 0 0
2
5.8993e-315 5.36716e-315
0
10 Polar Cap~
219 652 73 0 2 5
0 3 2
0
0 0 848 270
5 470uF
13 0 48 8
2 C3
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3723 0 0
2
5.8993e-315 5.3568e-315
0
9 I Source~
198 755 72 0 2 5
0 3 2
0
0 0 17264 0
5 4.0mA
20 0 55 8
3 Is3
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
6244 0 0
2
5.8993e-315 5.34643e-315
0
6 Diode~
219 623 45 0 2 5
0 4 3
0
0 0 848 0
6 1N4007
-21 -18 21 -10
2 D3
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6421 0 0
2
5.8993e-315 5.26354e-315
0
7 Ground~
168 610 102 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7743 0 0
2
5.8993e-315 0
0
7 Ground~
168 381 101 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9840 0 0
2
5.8993e-315 0
0
11 Signal Gen~
195 331 49 0 64 64
0 4 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1101004800 0 1103888384
0 814313567 814313567 981668463 1028443341 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 20 0 25.5 0 1e-09 1e-09 0.001 0.05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 0/25.5V
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
42 %D %1 %2 DC 0 PULSE(0 25.5 0 1n 1n 1m 50m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6910 0 0
2
5.8993e-315 5.26354e-315
0
6 Diode~
219 394 44 0 2 5
0 4 5
0
0 0 848 0
6 1N4007
-21 -18 21 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
449 0 0
2
5.8993e-315 0
0
7 Ground~
168 423 179 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8761 0 0
2
5.8993e-315 0
0
6 Diode~
219 423 135 0 2 5
0 2 6
0
0 0 848 90
6 1N4007
12 0 54 8
2 D2
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6748 0 0
2
5.8993e-315 0
0
9 I Source~
198 526 71 0 2 5
0 5 2
0
0 0 17264 0
5 4.0mA
20 0 55 8
3 Is2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
7393 0 0
2
5.8993e-315 5.3568e-315
0
10 Polar Cap~
219 423 72 0 2 5
0 5 2
0
0 0 848 270
5 470uF
13 0 48 8
2 C1
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7699 0 0
2
5.8993e-315 5.34643e-315
0
7 Ground~
168 422 101 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6638 0 0
2
5.8993e-315 5.32571e-315
0
7 Ground~
168 485 179 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4595 0 0
2
5.8993e-315 5.30499e-315
0
7 Ground~
168 526 101 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9395 0 0
2
5.8993e-315 5.26354e-315
0
9 Inductor~
219 485 145 0 2 5
0 6 2
0
0 0 848 270
3 1mH
6 -4 27 4
2 L1
10 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3303 0 0
2
5.8993e-315 0
0
7 Ground~
168 124 100 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4498 0 0
2
5.8993e-315 5.3568e-315
0
7 Ground~
168 83 100 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9728 0 0
2
5.8993e-315 5.34643e-315
0
7 Ground~
168 20 100 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
2
5.8993e-315 5.32571e-315
0
10 Polar Cap~
219 21 71 0 2 5
0 7 2
0
0 0 848 270
5 470uF
13 0 48 8
2 C2
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3978 0 0
2
5.8993e-315 5.30499e-315
0
9 I Source~
198 124 70 0 2 5
0 7 2
0
0 0 17264 0
5 4.0mA
20 0 55 8
3 Is1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
3494 0 0
2
5.8993e-315 5.26354e-315
0
4 .IC~
207 20 28 0 1 3
0 7
0
0 0 54096 0
3 25V
-11 -15 10 -7
4 CMD1
-13 -24 15 -16
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
3507 0 0
2
5.8993e-315 0
0
11 Resistor:A~
219 714 71 0 3 5
0 2 3 -1
0
0 0 880 90
3 330
7 3 28 11
2 R3
6 -8 20 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5151 0 0
2
5.8993e-315 5.39824e-315
0
11 Resistor:A~
219 485 70 0 2 5
0 6 5
0
0 0 880 90
3 330
7 3 28 11
2 R1
6 -8 20 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3701 0 0
2
5.8993e-315 5.36716e-315
0
11 Resistor:A~
219 83 69 0 3 5
0 2 7 -1
0
0 0 880 90
3 330
7 3 28 11
2 R2
6 -8 20 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8585 0 0
2
5.8993e-315 5.36716e-315
0
26
1 1 2 0 0 4096 0 25 1 0 0 2
714 89
714 94
1 0 3 0 0 4096 0 4 0 0 7 2
651 63
651 45
2 1 2 0 0 8320 0 0 7 0 0 3
591 55
610 55
610 96
1 0 4 0 0 12416 0 6 0 0 12 5
613 45
543 45
543 9
369 9
369 44
1 2 2 0 0 0 0 2 5 0 0 2
755 96
755 93
1 0 3 0 0 8192 0 5 0 0 7 3
755 51
755 45
714 45
2 2 3 0 0 8320 0 25 6 0 0 3
714 53
714 45
633 45
1 2 2 0 0 0 0 3 4 0 0 2
651 96
651 80
0 1 2 0 0 0 0 0 16 0 0 2
485 169
485 173
1 0 5 0 0 4096 0 14 0 0 19 2
422 62
422 44
2 1 2 0 0 0 0 9 8 0 0 3
362 54
381 54
381 95
1 1 4 0 0 0 0 10 9 0 0 2
384 44
362 44
1 1 2 0 0 0 0 12 11 0 0 2
423 145
423 173
2 0 6 0 0 8320 0 12 0 0 16 3
423 125
423 116
485 116
2 1 2 0 0 0 0 18 16 0 0 2
485 163
485 173
1 1 6 0 0 0 0 18 26 0 0 2
485 127
485 88
1 2 2 0 0 0 0 17 13 0 0 2
526 95
526 92
1 0 5 0 0 8192 0 13 0 0 19 3
526 50
526 44
485 44
2 2 5 0 0 8320 0 26 10 0 0 3
485 52
485 44
404 44
1 2 2 0 0 0 0 15 14 0 0 2
422 95
422 79
1 2 2 0 0 0 0 19 23 0 0 2
124 94
124 91
1 0 7 0 0 8192 0 23 0 0 23 3
124 49
124 43
83 43
2 0 7 0 0 8320 0 27 0 0 24 3
83 51
83 43
20 43
1 1 7 0 0 0 0 22 24 0 0 2
20 61
20 40
1 1 2 0 0 0 0 20 27 0 0 2
83 94
83 87
1 2 2 0 0 0 0 21 22 0 0 2
20 94
20 78
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.15 0.0001 0.0001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
