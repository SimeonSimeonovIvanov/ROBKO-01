CircuitMaker Text
5.6
Probes: 1
Is1_1
Transient Analysis
0 90 40 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 240 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.537855 0.500000
344 179 1190 520
9961490 0
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 119 97 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6966 0 0
2
41437.8 0
0
7 Ground~
168 78 97 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9796 0 0
2
41437.8 2
0
7 Ground~
168 15 97 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5952 0 0
2
41437.8 1
0
10 Polar Cap~
219 16 68 0 2 5
0 3 2
0
0 0 848 270
6 9400uF
10 0 52 8
2 C2
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3649 0 0
2
41437.8 0
0
9 I Source~
198 119 67 0 2 5
0 3 2
0
0 0 17264 0
5 300mA
13 0 48 8
3 Is1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 0 0 0 0
2 Is
3716 0 0
2
41437.8 0
0
4 .IC~
207 15 25 0 1 3
0 3
0
0 0 54096 0
3 15V
-11 -15 10 -7
4 CMD1
-13 -24 15 -16
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
4797 0 0
2
41437.8 0
0
11 Resistor:A~
219 78 66 0 3 5
0 2 3 -1
0
0 0 880 90
1 3
7 1 14 9
2 R2
6 -8 20 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4681 0 0
2
41437.8 3
0
6
1 2 2 0 0 4096 0 1 5 0 0 2
119 91
119 88
1 0 3 0 0 8192 0 5 0 0 3 3
119 46
119 40
78 40
2 0 3 0 0 8320 0 7 0 0 4 3
78 48
78 40
15 40
1 1 3 0 0 0 0 4 6 0 0 2
15 58
15 37
1 1 2 0 0 4096 0 2 7 0 0 2
78 91
78 84
1 2 2 0 0 4224 0 3 4 0 0 2
15 91
15 75
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.01 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
